/*Joshua Torres Morales A76478
  joshtm00@gmail.com*/

// MODE = 1 FIFO
// MODE = 0 LIFO

`include "ram.v"

module DUT #(parameter MODE=1'b1, parameter dat_width=32, parameter L=6, parameter DEPTH=64) 
(	input   [dat_width-1:0] Datain,
	input   Wren,
	input   Rden, 
	input   Wrclk,   
	input   Rdclk,   
	input   Rst,
	output  reg Full,
	output  reg Empty,
	output  reg [dat_width-1:0] Dataout
);   

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Internal Wires and Regs 
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

	wire [dat_width-1:0] data_ram;
	wire CLK;
  
	//Punteros de escritura y lectura, variable para contar datos en la memoria
	reg [L-1:0] adr_rd_i;
	reg [L-1:0] adr_wr_i;
	reg [L-1:0] status_cnt; 
  	
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 // Comb. Logic 
 //////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
   
	//Esto es para decidir cual reloj usar dependiedo del modo
	assign CLK = (MODE == 1'b1 )? Rdclk : Wrclk;
	//assign Dataout = data_ram;
  		
	
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Manejo del puntero de escritura
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	always @ (posedge Wrclk or posedge Rst) begin : WRITE_POINTER

		if (Rst) begin
			adr_wr_i <= 0;
		end 
		
		else if (Wrclk && Wren) begin
		
			if (adr_wr_i == DEPTH ) begin
				adr_wr_i <= adr_wr_i;
			end 
			
			else begin
				adr_wr_i <= adr_wr_i + 1;
			end
			
		end
		
		//In Stack Mode
		if((MODE==0) && Rden) begin
			
			if(adr_wr_i == 0) begin
				adr_wr_i <= adr_wr_i;
			end
			
			else begin		
				adr_wr_i <= adr_wr_i -1;
			end
		
		end
		
	end

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
//Manejo del puntero de lectura
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

	always @ (posedge CLK or posedge Rst) begin : READ_POINTER
	
		if (Rst) begin
			adr_rd_i <= 0;
		end 
		
		//In Queue Mode
		else if (Rden && (MODE == 1'b1) ) begin
			if (adr_rd_i == DEPTH ) begin
				adr_rd_i <= adr_rd_i;               
			end 
			
			else begin
				adr_rd_i <= adr_rd_i + 1;
         end    		
		end 
		
		//In Stack Mode, only one pointer is needed.		
		if(MODE == 1'b0) begin
			adr_rd_i <= adr_wr_i-1;
		end
		
	end
	
	
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Get the data from the RAM module	
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	

	always  @ (posedge CLK or posedge Rst ) begin : READ_DATA
		if (Rst ||!Rden ) begin
			Dataout <= 0;
		end else if (Rden) begin
			Dataout <= data_ram;
		end 
	end
	
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Status Counter
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	always @ (posedge CLK or posedge Rst) begin : STATUS_COUNTER
		
		//At Reset, the data structure is assumed empty.
		if (Rst) begin
			status_cnt <= 0;
		
		// If a Read command occurs, the Status Counter decreases by one.
		end else if (Rden &&  !(Wren) && (status_cnt  != 0) ) begin
			status_cnt <= status_cnt - 1;
			
		// If a Write command occurs:
		end else if (Wren &&  !(Rden) && (status_cnt  != DEPTH)) begin
			
			//If the Data Structure is full, the Status Counter stays the same.
			if (status_cnt == (DEPTH-1)) begin
				status_cnt <=status_cnt;
			
			//Else, the Status Counter increases by one  
			end else begin
				status_cnt <= status_cnt + 1;
			
			/*If both a Read and a Write commands occurs at the same time,
			the Status Counter increases and decreases by one, so no action is
			requiered.*/
			
			end
		end
	end 

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
//Syncronic Full and Empty signals.
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	always @ (posedge Wrclk or posedge Rst) begin: FULL_EMPTY
	
		if (Rst) begin
			Full  <= 0 ;
			Empty <= 1 ;

		end else if (status_cnt == (DEPTH-1)) begin
			Full  <= 1 ;
			Empty <= 0 ;
			
		end else if (status_cnt == 0) begin
			Full  <= 0 ;
			Empty <= 1 ;
		
		end else begin
			Full  <= 0 ;
			Empty <= 0 ;
		end
	end
	
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Ram instantiation, The ram is used as a data buffer.
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////		
	ram #(
		.mem_size(DEPTH),
		.adr_width(L),
		.dat_width(dat_width)
	) RAM(
			.dat_i(Datain), 
			.dat_o(data_ram), 
			.adr_wr_i(adr_wr_i), 
			.adr_rd_i(adr_rd_i), 
			.we_i(Wren), 
			.rde_i(Rden), 
			.clk(CLK)
			);
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
endmodule 
